`ifndef SNITCH_HWPE_SUBSYSTEM_SVH
`define SNITCH_HWPE_SUBSYSTEM_SVH


`define SNITCH_HWPE_SUBSYSTEM_BASE_ADDR 64'h00000000
`define SNITCH_HWPE_SUBSYSTEM_SIZE      64'h000000A0

`define SNITCH_HWPE_SUBSYSTEM_EVT_CLR_REG_ADDR   64'h00000094
`define SNITCH_HWPE_SUBSYSTEM_EVT_CLR_REG_OFFSET 64'h00000094

`define SNITCH_HWPE_SUBSYSTEM_MUX_SEL_REG_ADDR   64'h00000098
`define SNITCH_HWPE_SUBSYSTEM_MUX_SEL_REG_OFFSET 64'h00000098

`define SNITCH_HWPE_SUBSYSTEM_CLK_EN_REG_ADDR   64'h0000009C
`define SNITCH_HWPE_SUBSYSTEM_CLK_EN_REG_OFFSET 64'h0000009C


`endif /* SNITCH_HWPE_SUBSYSTEM_SVH */
